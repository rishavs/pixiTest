<?xml version="1.0" encoding="UTF-8"?>
<Batch version="1.0"><TaskList><Task type="ResizeTask" enabled="True"><Width units="0">64</Width><Height units="0">44</Height><DPI>-1</DPI><Filter>5</Filter><UseProportions>True</UseProportions></Task><Task type="ColorBalanceTask" enabled="True"><Red>19</Red><Green>0</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>40</Red><Green>0</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>59</Red><Green>0</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>80</Red><Green>0</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>98</Red><Green>0</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>2</Red><Green>19</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>2</Red><Green>38</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>2</Red><Green>59</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>2</Red><Green>79</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>2</Red><Green>97</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-18</Red><Green>1</Green><Blue>20</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-19</Red><Green>1</Green><Blue>38</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-39</Red><Green>-19</Green><Blue>18</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-59</Red><Green>-38</Green><Blue>19</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>20</Red><Green>-22</Green><Blue>38</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-18</Red><Green>-38</Green><Blue>39</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-19</Red><Green>0</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-39</Red><Green>-3</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-37</Red><Green>-55</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-35</Red><Green>-80</Green><Blue>0</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task><Task type="ColorBalanceTask" enabled="True"><Red>-98</Red><Green>-80</Green><Blue>-19</Blue></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><FileType></FileType><FilePath><![CDATA[C:\Users\rsharan\Desktop\test]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed></Task></TaskList></Batch>
